module page_bb(
    input wire clk_200,
    input wire clk_250,
    input wire clk_300, 
    input wire clk_350, 
    input wire clk_400, 
    input wire [48 : 0] din_leaf_bft2interface,
    output wire [48 : 0] dout_leaf_interface2bft,
    input wire resend,
    input wire reset_400,
    input wire ap_start
    );
    
endmodule
